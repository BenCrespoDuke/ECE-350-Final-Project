module servoController(clck,IR,DataA,DataB,Direction1,Direction2,Direction3,Direction4,Signals);

input clck;
input [31:0] DataA,DataB,IR;
output [1:0] Direction1,Direction2,Direction3,Direction4;
output [3:0] Signals;


endmodule