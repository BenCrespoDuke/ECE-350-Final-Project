module MoveMem(
    IR_In, DirIn, SpeedIn, Shift,clck,reset
);



register dir1(data_In, data_Out, clk,en,clr);
register speed1(data_In, data_Out, clk,en,clr);
register dir1(data_In, data_Out, clk,en,clr);
register speed1(data_In, data_Out, clk,en,clr);
register dir1(data_In, data_Out, clk,en,clr);
register speed1(data_In, data_Out, clk,en,clr);
register dir1(data_In, data_Out, clk,en,clr);
register speed1(data_In, data_Out, clk,en,clr);
endmodule