module LeftShifter(dataA,shiftAm,out);
     input[31:0] dataA;
     input [4:0] shiftAm;
     output[31:0] out;
     wire [31:0] w1,w2,w3,w4,w5,w6,w7,w8,w9;
     and sn161(w1[0],0,dataA[0]);
     and sn162(w1[1],0,dataA[0]);
     and sn163(w1[2],0,dataA[0]);
     and sn164(w1[3],0,dataA[0]);
     and sn165(w1[4],0,dataA[0]);
     and sn166(w1[5],0,dataA[0]);
     and sn167(w1[6],0,dataA[0]);
     and sn168(w1[7],0,dataA[0]);
     and sn169(w1[8],0,dataA[0]);
     and sn1610(w1[9],0,dataA[0]);
     and sn1611(w1[10],0,dataA[0]);
     and sn1612(w1[11],0,dataA[0]);
     and sn1613(w1[12],0,dataA[0]);
     and sn1614(w1[13],0,dataA[0]);
     and sn1615(w1[14],0,dataA[0]);
     and sn1616(w1[15],0,dataA[0]);

     and s161(w1[16],1,dataA[0]);
     and s162(w1[17],1,dataA[1]);
     and s163(w1[18],1,dataA[2]);
     and s164(w1[19],1,dataA[3]);
     and s165(w1[20],1,dataA[4]);
     and s166(w1[21],1,dataA[5]);
     and s167(w1[22],1,dataA[6]);
     and s168(w1[23],1,dataA[7]);
     and s169(w1[24],1,dataA[8]);
     and s1610(w1[25],1,dataA[9]);
     and s1611(w1[26],1,dataA[10]);
     and s1612(w1[27],1,dataA[11]);
     and s1613(w1[28],1,dataA[12]);
     and s1614(w1[29],1,dataA[13]);
     and s1615(w1[30],1,dataA[14]);
     and s1616(w1[31],1,dataA[15]);
     
     mux_2 is16(w2,shiftAm[4],dataA,w1);

     and sn81(w3[0],0,w2[0]);
     and sn82(w3[1],0,w2[0]);
     and sn83(w3[2],0,w2[0]);
     and sn84(w3[3],0,w2[0]);
     and sn85(w3[4],0,w2[0]);
     and sn86(w3[5],0,w2[0]);
     and sn87(w3[6],0,w2[0]);
     and sn88(w3[7],0,w2[0]);
     and sn89(w3[8],1,w2[0]);
     and sn810(w3[9],1,w2[1]);
     and sn811(w3[10],1,w2[2]);
     and sn812(w3[11],1,w2[3]);
     and sn813(w3[12],1,w2[4]);
     and sn814(w3[13],1,w2[5]);
     and sn815(w3[14],1,w2[6]);
     and sn816(w3[15],1,w2[7]);

     and s81(w3[16],1,w2[8]);
     and s82(w3[17],1,w2[9]);
     and s83(w3[18],1,w2[10]);
     and s84(w3[19],1,w2[11]);
     and s85(w3[20],1,w2[12]);
     and s86(w3[21],1,w2[13]);
     and s87(w3[22],1,w2[14]);
     and s88(w3[23],1,w2[15]);
     and s89(w3[24],1,w2[16]);
     and s810(w3[25],1,w2[17]);
     and s811(w3[26],1,w2[18]);
     and s812(w3[27],1,w2[19]);
     and s813(w3[28],1,w2[20]);
     and s814(w3[29],1,w2[21]);
     and s815(w3[30],1,w2[22]);
     and s816(w3[31],1,w2[23]);

     mux_2 is8(w4,shiftAm[3],w2,w3);

     and sn41(w5[0],0,w4[0]);
     and sn42(w5[1],0,w4[0]);
     and sn43(w5[2],0,w4[0]);
     and sn44(w5[3],0,w4[0]);
     and sn45(w5[4],1,w4[0]);
     and sn46(w5[5],1,w4[1]);
     and sn47(w5[6],1,w4[2]);
     and sn48(w5[7],1,w4[3]);
     and sn49(w5[8],1,w4[4]);
     and sn410(w5[9],1,w4[5]);
     and sn411(w5[10],1,w4[6]);
     and sn412(w5[11],1,w4[7]);
     and sn413(w5[12],1,w4[8]);
     and sn414(w5[13],1,w4[9]);
     and sn415(w5[14],1,w4[10]);
     and sn416(w5[15],1,w4[11]);

     and s41(w5[16],1,w4[12]);
     and s42(w5[17],1,w4[13]);
     and s43(w5[18],1,w4[14]);
     and s44(w5[19],1,w4[15]);
     and s45(w5[20],1,w4[16]);
     and s46(w5[21],1,w4[17]);
     and s47(w5[22],1,w4[18]);
     and s48(w5[23],1,w4[19]);
     and s49(w5[24],1,w4[20]);
     and s410(w5[25],1,w4[21]);
     and s411(w5[26],1,w4[22]);
     and s412(w5[27],1,w4[23]);
     and s413(w5[28],1,w4[24]);
     and s414(w5[29],1,w4[25]);
     and s415(w5[30],1,w4[26]);
     and s416(w5[31],1,w4[27]);

     mux_2 is4(w6,shiftAm[2],w4,w5);

     and sn21(w7[0],0,w6[0]);
     and sn22(w7[1],0,w6[0]);
     and sn23(w7[2],1,w6[0]);
     and sn24(w7[3],1,w6[1]);
     and sn25(w7[4],1,w6[2]);
     and sn26(w7[5],1,w6[3]);
     and sn27(w7[6],1,w6[4]);
     and sn28(w7[7],1,w6[5]);
     and sn29(w7[8],1,w6[6]);
     and sn210(w7[9],1,w6[7]);
     and sn211(w7[10],1,w6[8]);
     and sn212(w7[11],1,w6[9]);
     and sn213(w7[12],1,w6[10]);
     and sn214(w7[13],1,w6[11]);
     and sn215(w7[14],1,w6[12]);
     and sn216(w7[15],1,w6[13]);

     and s21(w7[16],1,w6[14]);
     and s22(w7[17],1,w6[15]);
     and s23(w7[18],1,w6[16]);
     and s24(w7[19],1,w6[17]);
     and s25(w7[20],1,w6[18]);
     and s26(w7[21],1,w6[19]);
     and s27(w7[22],1,w6[20]);
     and s28(w7[23],1,w6[21]);
     and s29(w7[24],1,w6[22]);
     and s210(w7[25],1,w6[23]);
     and s211(w7[26],1,w6[24]);
     and s212(w7[27],1,w6[25]);
     and s213(w7[28],1,w6[26]);
     and s214(w7[29],1,w6[27]);
     and s215(w7[30],1,w6[28]);
     and s216(w7[31],1,w6[29]);

    mux_2 is2(w8,shiftAm[1],w6,w7);

    and sn11(w9[0],0,w8[0]);
     and sn12(w9[1],1,w8[0]);
     and sn13(w9[2],1,w8[1]);
     and sn14(w9[3],1,w8[2]);
     and sn15(w9[4],1,w8[3]);
     and sn16(w9[5],1,w8[4]);
     and sn17(w9[6],1,w8[5]);
     and sn18(w9[7],1,w8[6]);
     and sn19(w9[8],1,w8[7]);
     and sn110(w9[9],1,w8[8]);
     and sn111(w9[10],1,w8[9]);
     and sn112(w9[11],1,w8[10]);
     and sn113(w9[12],1,w8[11]);
     and sn114(w9[13],1,w8[12]);
     and sn115(w9[14],1,w8[13]);
     and sn116(w9[15],1,w8[14]);

     and s11(w9[16],1,w8[15]);
     and s12(w9[17],1,w8[16]);
     and s13(w9[18],1,w8[17]);
     and s14(w9[19],1,w8[18]);
     and s15(w9[20],1,w8[19]);
     and s16(w9[21],1,w8[20]);
     and s17(w9[22],1,w8[21]);
     and s18(w9[23],1,w8[22]);
     and s19(w9[24],1,w8[23]);
     and s110(w9[25],1,w8[24]);
     and s111(w9[26],1,w8[25]);
     and s112(w9[27],1,w8[26]);
     and s113(w9[28],1,w8[27]);
     and s114(w9[29],1,w8[28]);
     and s115(w9[30],1,w8[29]);
     and s116(w9[31],1,w8[30]);

     mux_2 is1(out,shiftAm[0],w8,w9);

endmodule